// ----------------------------------------------------------------------------
//
// ----------------------------------------------------------------------------
// FILE NAME      : sl_core_inc.sv
// PROJECT        : Selen
// AUTHOR         : Grigoriy Zhikharev
// AUTHOR'S EMAIL : gregory.zhiharev@gmail.com
// ----------------------------------------------------------------------------
// DESCRIPTION    :
// ----------------------------------------------------------------------------

`ifndef INC_SL_CORE_INC
`define INC_SL_CORE_INC

`include "core/sl_core_if.sv"
`include "core/sl_core_typedefs.sv"
`include "core/sl_core_bus_item.sv"
`include "core/sl_core_agent_cfg.sv"
`include "core/sl_core_monitor.sv"
`include "core/sl_core_sequencer.sv"
`include "core/sl_core_slave_driver.sv"
`include "core/sl_core_slave_agent.sv"
`include "core/sl_core_master_driver.sv"
`include "core/sl_core_master_agent.sv"
`include "core/sl_core_seq_lib.sv"

`endif
