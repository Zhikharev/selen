// ----------------------------------------------------------------------------
//
// ----------------------------------------------------------------------------
// FILE NAME      : sl_wb_inc.sv
// PROJECT        : Selen
// AUTHOR         : Maksim Kobzar
// AUTHOR'S EMAIL : maksim.s.kobzar@gmail.com
// ----------------------------------------------------------------------------
// DESCRIPTION    :
// ----------------------------------------------------------------------------

`ifndef INC_SL_WB_INC
`define INC_SL_WB_INC

`include "wishbone/sl_wb_defines.sv"
`include "wishbone/sl_wb_interface.sv"
`include "wishbone/sl_wb_agent_cfg.sv"
`include "wishbone/sl_wb_bus_item.sv"
`include "wishbone/sl_wb_monitor.sv"
`include "wishbone/sl_wb_sequencer.sv"
`include "wishbone/sl_wb_slave_driver.sv"
`include "wishbone/sl_wb_slave_agent.sv"

`endif
