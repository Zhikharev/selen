
module io_top();

endmodule