`define WB_DATA_WIDTH 	32
`define WB_ADDR_WIDTH 	32
`define WB_BE_WIDTH   	(`WB_DATA_WIDTH/8)