
$GIT_HOME/rtl/lib/fifo.v
$GIT_HOME/rtl/lib/sram_sp.v
$GIT_HOME/rtl/lib/sram_dp.v
$GIT_HOME/rtl/l1_cache/l1_defines.sv
$GIT_HOME/rtl/l1_cache/l1_lrum.sv
$GIT_HOME/rtl/l1_cache/l1_ld_mem.sv
$GIT_HOME/rtl/l1_cache/l1_dm_mem.sv
$GIT_HOME/rtl/l1_cache/l1_mau.sv
$GIT_HOME/rtl/l1_cache/l1i_top.sv
$GIT_HOME/rtl/l1_cache/l1d_top.sv
