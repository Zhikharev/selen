// ----------------------------------------------------------------------------
//
// ----------------------------------------------------------------------------
// FILE NAME      : selen_tb_top.sv
// PROJECT        : Selen
// AUTHOR         : Grigoriy Zhikharev
// AUTHOR'S EMAIL : gregory.zhiharev@gmail.com
// ----------------------------------------------------------------------------
// DESCRIPTION    :
// ----------------------------------------------------------------------------

`ifndef INC_SELEN_TB_TOP
`define INC_SELEN_TB_TOP

`ifndef CLK_HALF_TIME
`define CLK_HALF_TIME 16ns
`endif

`define CORE_PATH selen_top.cpu_cluster.core

module selen_tb_top ();

	logic clk;
	logic rst;

	wire gpio_pin_o;
	wire gpio_pin_en;
	wire gpio_pin_i;

	tri gpio_bus;

	assign gpio_pin_i = gpio_bus;
	assign gpio_bus = (gpio_pin_en) ? gpio_pin_o : 1'bZ;

  wire   spi_ss;
  wire   spi_sclk;
  wire   spi_mosi;
  wire   spi_miso;

	initial begin
		$display("CLK_HALF_TIME=%0d", `CLK_HALF_TIME);
		clk = 0;
		forever #`CLK_HALF_TIME clk = !clk;
	end

	initial	 begin
		rst = 1;
		repeat(5) @(posedge clk);
		rst = 0;
	end

	initial begin
		forever begin
			@(negedge clk);
			if(`CORE_PATH.d_req_val && `CORE_PATH.d_req_cop inside {0, 3}) begin
				do begin
					@(negedge clk);
				end
				while(!`CORE_PATH.d_req_ack);
				if(!$test$plusargs("NO_FATAL_ON_X")) begin
					if($isunknown(`CORE_PATH.d_ack_rdata)) #100 $fatal("Found X on d_ack_rdata after read operation");
				end
			end
		end
	end

	initial begin
		forever begin
			if(~rst) begin
				@(negedge clk);
				if(selen_top.cpu_cluster.core.i_req_val) begin
					string str;
					rv32_transaction item = new("item");
					str = {$sformatf("[INSTR] ADDR=%32h ", selen_top.cpu_cluster.core.i_req_addr)};
					while(!selen_top.cpu_cluster.core.i_req_ack) @(negedge clk);
					forever begin
						item.decode(selen_top.cpu_cluster.core.i_ack_rdata);
						str = {str, $sformatf("DATA=%32h ",selen_top.cpu_cluster.core.i_ack_rdata)};
						str = {str, item.sprint()};
						if($test$plusargs("INSTR_TRACE")) $display("%0s (%0t)", str, $time());
						str = {$sformatf("[INSTR] ADDR=%32h ", selen_top.cpu_cluster.core.i_req_addr)};
						do begin @(negedge clk);
						end
						while(!selen_top.cpu_cluster.core.i_req_ack);
					end
				end
			end
			else @(negedge clk);
		end
	end

	selen_top selen_top
	(
		.clk 					(clk),
		.rst_n 				(!rst),
		.gpio_pin0_o 	(),
		.gpio_pin0_en (),
		.gpio_pin0_i 	(1'b1),
		.gpio_pin1_o 	(gpio_pin_o),
		.gpio_pin1_en (gpio_pin_en),
		.gpio_pin1_i 	(gpio_pin_i),
  	.spi_ss_o 		(spi_ss),
  	.spi_sclk_o 	(spi_sclk),
  	.spi_mosi_o 	(spi_mosi),
  	.spi_miso_i 	(spi_miso)
	);

 	N25Qxxx spi_flash
 	(
 		.S  				(spi_ss),
 		.C_  				(spi_sclk),
 		.HOLD_DQ3 	(1'b1),
 		.DQ0 				(spi_mosi),
 		.DQ1 				(spi_miso),
 		.Vcc 				('d3000),
 		.Vpp_W_DQ2 	(1'b1)
 	);

	initial begin
		$display("%0t TEST START", $time());
		wait(selen_top.cpu_cluster.core.d_req_val && selen_top.cpu_cluster.core.d_req_addr == 32'hffff_fff0);
		$display("%0t TEST FINISHED", $time());
		$finish();
	end

  initial $timeformat(-9, 1, "ns", 4);

  `ifdef WAVES_FSDB
  initial begin
    $fsdbDumpfile("sl_tb_top");
    $fsdbDumpvars;
  end
  `elsif WAVES_VCD
  initial begin
     $dumpvars;
  end
  `elsif WAVES
  initial begin
    $vcdpluson;
  end
  `endif

  // -----------------------------------------
  // ROM IMAGE
  // -----------------------------------------
  initial $readmemh("rom_image.v", selen_top.wb_rom_5kB.rom.rom);
  initial $readmemh("ram_image.v", selen_top.wb_ram_256kB.ram.ram);

endmodule

`endif
