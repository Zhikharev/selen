// ----------------------------------------------------------------------------
//
// ----------------------------------------------------------------------------
// FILE NAME      : wb_inc.sv
// PROJECT        : Selen
// AUTHOR         : Maksim Kobzar
// AUTHOR'S EMAIL : maksim.s.kobzar@gmail.com
// ----------------------------------------------------------------------------
// DESCRIPTION    :
// ----------------------------------------------------------------------------

`ifndef INC_WB_INC
`define INC_WB_INC

`include "wishbone/wb_if.sv"
`include "wishbone/wb_agent_cfg.sv"
`include "wishbone/wb_item.sv"
`include "wishbone/wb_monitor.sv"
`include "wishbone/wb_sequencer.sv"
`include "wishbone/wb_slave_driver.sv"
`include "wishbone/wb_slave_agent.sv"

`endif
