module wb_data(
	input[31:0] data_in,
	input[31:0] addr2mem,
	output[31:0] data_out,
	input sw,
	input lw,
	input clk,
	input rst,
	output stb,
	input ack,
	input stall
);


endmodule
