// ----------------------------------------------------------------------------
// 
// ----------------------------------------------------------------------------
// FILE NAME      : cpu_assembled.sv
// PROJECT        : Selen
// AUTHOR         : 
// AUTHOR'S EMAIL : 
// ----------------------------------------------------------------------------
// DESCRIPTION    : 
// ----------------------------------------------------------------------------

`ifndef INC_CPU_ASSEMBLED
`define INC_CPU_ASSEMBLED

module cpu_assembled (
	input 				clk,
	input 				rst,
	wishbone_if 	wbi_intf,
	wishbone_if 	wbd_intf
);

	// Instantiate CPU DUT here

endmodule

`endif