// ----------------------------------------------------------------------------
// 
// ----------------------------------------------------------------------------
// FILE NAME      : wishbone_if.sv
// PROJECT        : Selen
// AUTHOR         : 
// AUTHOR'S EMAIL : 
// ----------------------------------------------------------------------------
// DESCRIPTION    : 
// ----------------------------------------------------------------------------

`ifndef INC_WISHBONE_IF
`define INC_WISHBONE_IF

interface wishbone_if (input logic clk, input logic rst);
endinterface

`endif