`include "uvm_pkg.sv"
`include "uvm_macros.svh"

`include "testbench/l1_rtl_inc.sv"

`include "wb_if.sv"
`include "sl_core_if.sv"

import uvm_pkg::*;

`include "uvm/uvm.inc.sv"
`include "testbench/l1_assembled.sv"
`include "testbench/l1_tb_top.sv"
