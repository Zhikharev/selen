// ----------------------------------------------------------------------------
// 
// ----------------------------------------------------------------------------
// FILE NAME      : core_assembled.sv
// PROJECT        : Selen
// AUTHOR         : 
// AUTHOR'S EMAIL : 
// ----------------------------------------------------------------------------
// DESCRIPTION    : 
// ----------------------------------------------------------------------------

`ifndef INC_CORE_ASSEMBLED
`define INC_CORE_ASSEMBLED


module core_assembled (
	input 				clk,
	input 				rst,
	core_if 			i_intf,
	core_if 			d_intf
);


	// Instantiate CPU DUT here


endmodule

`endif
