`ifndef INC_RST_IFC_MODEL_INC
`define INC_RST_IFC_MODEL_INC

`include "rst_ifc/rst_model_driver.sv"

`endif