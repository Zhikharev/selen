// ----------------------------------------------------------------------------
// 
// ----------------------------------------------------------------------------
// FILE NAME      : cpu_assembled.sv
// PROJECT        : Selen
// AUTHOR         : 
// AUTHOR'S EMAIL : 
// ----------------------------------------------------------------------------
// DESCRIPTION    : 
// ----------------------------------------------------------------------------

`ifndef INC_CPU_ASSEMBLED
`define INC_CPU_ASSEMBLED

module cpu_assembled (
	input 				clk,
	input 				rst,
	wishborne_if 	wbi_intf,
	wishborne_if 	wbd_intf
);

	// Instantiate CPU DUT here

endmodule

`endif