`ifndef INC_RST_IFC_INC
`define INC_RST_IFC_INC

`include "rst_ifc/rst_interface.sv"
`include "rst_ifc/rst_transfer_item.sv"
`include "rst_ifc/rst_driver.sv"
`include "rst_ifc/rst_monitor.sv"
`include "rst_ifc/rst_agent.sv"
`include "rst_ifc/rst_base_seq.sv"

`endif