// ----------------------------------------------------------------------------
//
// ----------------------------------------------------------------------------
// FILE NAME      : sl_core_sequencer.sv
// PROJECT        : Selen
// AUTHOR         :
// AUTHOR'S EMAIL :
// ----------------------------------------------------------------------------
// DESCRIPTION    :
// ----------------------------------------------------------------------------

`ifndef INC_SL_CORE_SEQUENCER
`define INC_SL_CORE_SEQUENCER

typedef uvm_sequencer#(sl_core_bus_item) sl_core_sequencer;

`endif
