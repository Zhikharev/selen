typedef enum int {
	ADD
} r32v_opcode;