`define R_OPCODE 7'b0110011
`define I_R_OPCODE 7'b0010011
`define LUI_OPCODE 7'b0110111
`define AUIPC_OPCODE 7'b0010111
`define SB_OPCODE 7'b1100011
`define UJ_OPCODE 7'b1101111
`define JALR_OPCODE 7'b1100111
`define LD_OPCODE 7'b0000011
`define ST_OPCODE 7'b0100011

`define FNCT7_1 7'b0
`define FNCT7_2 7'b0100000

`define ADD 3'b000
`define SLT 3'b010
`define SLTU 3'b011
`define AND	3'b111
`define OR 3'b110
`define XOR 3'b100
`define SLL 3'b001
`define SRL 3'b101
`define SUB	3'b000
`define SRA 3'b101
`define AM	3'b010

`define ADDI 3'b000
`define SLTI 3'b010
`define SLTUI 3'b011
`define ANDI 3'b111
`define ORI 3'b110
`define XORI 3'b100
`define SLLI 3'b001
`define SRLI 3'b101
`define SRAI 3'b101

`define BEQ 3'b000
`define BNE 3'b001
`define BLT 3'b100
`define BLTU 3'b110
`define BGE 3'b101
`define BGEU 3'b111

`define JALR 3'b000
`define LH 3'b001
`define LW 3'b010
`define LHU 3'b101
`define LBU 3'b100
`define  LB 3'b000 

`define SW 3'b010
`define SH 3'b001
`define SB 3'b000

