`ifndef UVM_INC
`define UVM_INC

`include "uvm_pkg.sv"
`include "uvm_macros.svh"

import uvm_pkg::*;

// Common
`include "smart_report_server.sv"
`include "core/sl_core_inc.sv"

`endif