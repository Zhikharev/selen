typedef enum int {
	ADD
} rv32_opcode;